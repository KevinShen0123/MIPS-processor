module sx(result, immed);
input[16:0] immed
output [31:0] data_result
wire isNotEqual,isLessThan,overflow
alu(immed, immed, 5'b00101, 5'b10000, data_result, isNotEqual, isLessThan, overflow);




endmodule